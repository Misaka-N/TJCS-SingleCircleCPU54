`timescale 1ns / 1ps
module PC(                      //ָ���ַ�Ĵ���
    input  pc_clk,              //PC�Ĵ�����ʱ���źţ�д��Ϊͬ����ʱ���½�����Ч������ȡΪ�첽
    input  pc_ena,              //ʹ�ܶ��źţ��ߵ�ƽ��Ч
    input  rst,                 //��λ�źţ��ߵ�ƽ��Ч
    input  [31:0] pc_addr_in,   //��������PC�Ĵ�����ָ���ַ��Ҳ������һ��Ҫִ�е�ָ��
    output [31:0] pc_addr_out   //���δ�PC�Ĵ����д�����ָ���ַ��Ҳ���ǵ�ǰ��Ҫִ�е�ָ��
    );
/* �ڲ��ñ��� */
reg [31:0] pc_reg = 32'h00400000;//��ʼλ����32'h00400000����˸���ֵҲ�����

/* ��ֵ���첽��ȡ */
assign pc_addr_out = pc_ena ? pc_reg : 32'hz;   //ֻҪʹ�ܶ�Ϊ�ߵ�ƽ������PC�Ĵ���������ʱ���Զ�ȡ����

/* �����������첽д������� */
always @(negedge pc_clk or posedge rst)   //��λ�ź������ػ�ʱ���½�����Ч
begin
    if(rst && pc_ena)           //��λ�źŸߵ�ƽ����λ��ȫ����0������������д������ena����ֻ�����üĴ����Ѻ������գ����Ӵ�����ʱ���ԣ�Ϊ�����ݰ�ȫ���ǣ��������ǰ�ߣ���ֹ�Ĵ������ݱ���������գ�
        pc_reg <= 32'h00400000; //ע����ʼλ��ʱ32'h00400000
    else if(pc_ena)             //��ִ�е�����˵��clk�����½��أ�ֻҪʹ�ܶ�Ϊ�ߵ�ƽ�Ϳ��޸�PC��ֵ
        pc_reg <= pc_addr_in;

end

endmodule
